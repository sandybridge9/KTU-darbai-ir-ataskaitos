------------------------------------- 

--KTU 2015

--Informatikos fakultetas
--Kompiuteriu katedra
--Kompiuteriu Architektura [P175B125] 
--Kazimieras Bagdonas 

--v1.0

------------------------------------- 
--KTU 2016 

--ditto

--v1.01
--panaikinta "save" mikrokomanda registrams, sutrumpinta ROM eilute nuo 75 iki 69 bitu, nesuderinama su V1.0   

------------------------------------- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is 
	port (
		RST_ROM : in std_logic;
		ROM_CMD : in std_logic_vector(7 downto 0);  
		ROM_Dout : out std_logic_vector(1 to 69)
		);
end ROM ;

architecture rtl of ROM is
	
	type memory is array (0 to 255) of std_logic_vector(1 to 69) ; 
	
	constant ROM_CMDln : memory := (  
--                    1         2         3         4         5         6            Dvi komentaro eilutes duoda bitu numerius   
--           123456789012345678901234567890123456789012345678901234567890123456789    (nuo 1 iki 69)
	0=> "010000000000000100000000000000000000000000000000000000000000000000000",  --skaitom B
	1=> "000100000000000000000010000000000000000000000000000000000000000000000",  --C = B
	2=> "000000000000000000000000000000000000000000000000000000000010000000000",  --reset A
	3=> "101100000010100000000000000000000000000000000000000000000000000000000",  --LS = 6 (C Low = 1?)
	4=> "000100001000000000000000000000000000000000000000001000000000000000000",  --A = A + B
	5=> "000000000000000010000000100000000000000000000000000000000000000000001",  --LL1(B) LR1(C) CNT--
	6=> "111010000001100000000000000000000000000000000000000000000000000000000",  --LS = 13 (CNT = 0)
	7=> "001000000000000000000000000000000000000000000000000000000000000000010",  --rezultatas
	8=> "001000000000000000000000000000000000000000000000000000000000000000010",  --rezultatas
	9=> "010000000000000000000000000001000000000000000000000000000000000000000",  --D = Din
	10=> "001000000000000000000000000000000000100000000000000000000000000000000",  --E = A
	11=> "000000000000000000000000000000000000000000000000000000000010000000000",  --reset A
	12=> "000001001000000000000000000000000000000000000000000000000000000000000",  --A = D
	13=> "000000101000000000000000000000000000000000000000001000000000000000000",  --A = A + E
	14=> "001000000000000000000000000000000000000000000000000000000000000000010",  --rezultatas
	15=> "001000000000000000000000000000000000000000000000000000000000000000010",  --rezultatas


	
	others => (others => '0') );   
	
	
	
begin
	process (RST_ROM, ROM_CMD) 
		
	begin
		if RST_ROM'event and RST_ROM = '1' then 
			ROM_Dout <= ROM_CMDln(0);
		elsif ROM_CMD'event then
			ROM_Dout <= ROM_CMDln(to_integer(unsigned(ROM_CMD))); 
		end if;
		
	end process;
	
end rtl;